** Profile: "CC_2-Current sweep"  [ d:\projekty\power_supply\pcb_design\simulations\summing node-pspicefiles\cc_2\current sweep.sim ] 

** Creating circuit file "Current sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\David\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V10 3.3V 0V 0.1V 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\CC_2.net" 


.END
