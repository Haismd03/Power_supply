** Profile: "CC-Voltage sweep, I set"  [ D:\Projekty\Power_supply\PCB_design\Simulations\summing node-pspicefiles\cc\voltage sweep, i set.sim ] 

** Creating circuit file "Voltage sweep, I set.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\David\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM V_set 0 3.3 10m 
.STEP PARAM I_set LIST 3.0, 2.2, 1.2, 0.2, 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\CC.net" 


.END
