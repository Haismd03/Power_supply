** Profile: "CC_2-R_out sweep"  [ d:\projekty\power_supply\pcb_design\simulations\summing node-PSpiceFiles\CC_2\R_out sweep.sim ] 

** Creating circuit file "R_out sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\David\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM R_out 10 100m 100m 
.STEP PARAM I_node LIST 3, 2, 1, 0.5 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\CC_2.net" 


.END
