** Profile: "CC-Resistive sweep, I set"  [ D:\Projekty\Power_supply\PCB_design\Simulations\summing node-pspicefiles\cc\resistive sweep, i set.sim ] 

** Creating circuit file "Resistive sweep, I set.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\David\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM R_out 10 0.1 0.1 
.STEP LIN PARAM I_set 0.8 1.8 0.5 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\CC.net" 


.END
