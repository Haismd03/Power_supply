** Profile: "CC-Resistive sweep"  [ d:\projekty\power_supply\pcb_design\simulations\summing node-pspicefiles\cc\resistive sweep.sim ] 

** Creating circuit file "Resistive sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\David\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM R_out 10 0.1 0.01 
.STEP LIN PARAM V_node 1 3.2 0.5 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\CC.net" 


.END
