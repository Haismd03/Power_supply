** Profile: "summing node-V set, R sweep"  [ d:\projekty\power_supply\pcb_design\simulations\summing node-PSpiceFiles\summing node\V set, R sweep.sim ] 

** Creating circuit file "V set, R sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\David\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM V_node 3.3V 0V 0.1V 
.STEP LIN PARAM R_sweep 10 0.1 0.1 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\summing node.net" 


.END
