** Profile: "CC-Voltage sweep, low I"  [ d:\projekty\power_supply\pcb_design\simulations\summing node-pspicefiles\cc\voltage sweep, low i.sim ] 

** Creating circuit file "Voltage sweep, low I.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\David\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM V_set 3.3 0 0.05 
+ PARAM R_out LIST 1k 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\CC.net" 


.END
